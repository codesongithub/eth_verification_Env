class eth_cfg;
	static mailbox gen2bfm_mb= new();
	static mailbox bfm2gen_mb=new();
endclass
